module main

struct Settings {
	mut:
		location string
		api_key string
}