// Settings file for holding the City ID and API Key

module main

struct Settings {
	mut:
		location string
		api_key string
}