module main

struct VVeatherSettings {
	mut:
		location string
		api_key string
}